module uart_rx #(
    parameter
    /*
     You can specify the following three parameters.
     1. DATA_WIDTH : width of data that is transmited by this module
     2. BAUD_RATE  : baud rate of output uart signal
     3. CLK_FREQ   : freqency of input clock signal




    */
    DATA_WIDTH = 8,
    BAUD_RATE = 9600,
    CLK_FREQ = 12_000_000,

    localparam LB_DATA_WIDTH    = $clog2(DATA_WIDTH),
               PULSE_WIDTH      = CLK_FREQ / BAUD_RATE,
               LB_PULSE_WIDTH   = $clog2(PULSE_WIDTH),
               HALF_PULSE_WIDTH = PULSE_WIDTH / 2
) (
    input  logic                  sig,
    input  logic                  ready,
    output logic [DATA_WIDTH-1:0] data,
    output logic                  valid,
    input  logic                  clk,
    input  logic                  rstn
);

  //-----------------------------------------------------------------------------
  // noise removing filter



  function majority5(input [4:0] val);
    case (val)
      5'b00000: majority5 = 0;
      5'b00001: majority5 = 0;
      5'b00010: majority5 = 0;
      5'b00100: majority5 = 0;
      5'b01000: majority5 = 0;
      5'b10000: majority5 = 0;
      5'b00011: majority5 = 0;
      5'b00101: majority5 = 0;
      5'b01001: majority5 = 0;
      5'b10001: majority5 = 0;
      5'b00110: majority5 = 0;
      5'b01010: majority5 = 0;
      5'b10010: majority5 = 0;
      5'b01100: majority5 = 0;
      5'b10100: majority5 = 0;
      5'b11000: majority5 = 0;
      default:  majority5 = 1;
    endcase
  endfunction

  //-----------------------------------------------------------------------------
  // description about input signal



  logic [1:0] sampling_cnt;
  logic [4:0] sig_q;
  logic       sig_r;

  always_ff @(posedge clk) begin
    if (!rstn) begin
      sampling_cnt <= 0;
      sig_q        <= 5'b11111;
      sig_r        <= 1;
    end else begin
      // connect to deserializer after removing noise



      if (sampling_cnt == 0) begin
        sig_q <= {sig, sig_q[4:1]};
      end

      sig_r        <= majority5(sig_q);
      sampling_cnt <= sampling_cnt + 1;
    end
  end

  //----------------------------------------------------------------
  // description about receive UART signal



  typedef enum logic [1:0] {
    STT_DATA,
    STT_STOP,
    STT_WAIT
  } statetype;

  statetype                    state;

  logic     [  DATA_WIDTH-1:0] data_tmp_r;
  logic     [ LB_DATA_WIDTH:0] data_cnt;
  logic     [LB_PULSE_WIDTH:0] clk_cnt;
  logic                        rx_done;

  always_ff @(posedge clk) begin
    if (!rstn) begin
      state      <= STT_WAIT;
      data_tmp_r <= 0;
      data_cnt   <= 0;
      clk_cnt    <= 0;
    end else begin

      //-----------------------------------------------------------------------------
      // 3-state FSM



      case (state)

        //-----------------------------------------------------------------------------
        // state      : STT_DATA
        // behavior   : deserialize and recieve data
        // next state : when all data have recieved -> STT_STOP



        STT_DATA: begin
          if (0 < clk_cnt) begin
            clk_cnt <= clk_cnt - 1;
          end else begin
            data_tmp_r <= {sig_r, data_tmp_r[DATA_WIDTH-1:1]};
            clk_cnt    <= PULSE_WIDTH;

            if (data_cnt == DATA_WIDTH - 1) begin
              state <= STT_STOP;
            end else begin
              data_cnt <= data_cnt + 1;
            end
          end
        end

        //-----------------------------------------------------------------------------
        // state      : STT_STOP
        // behavior   : watch stop bit
        // next state : STT_WAIT



        STT_STOP: begin
          if (0 < clk_cnt) begin
            clk_cnt <= clk_cnt - 1;
          end else if (sig_r) begin
            state <= STT_WAIT;
          end
        end

        //-----------------------------------------------------------------------------
        // state      : STT_WAIT
        // behavior   : watch start bit
        // next state : when start bit is observed -> STT_DATA



        STT_WAIT: begin
          if (sig_r == 0) begin
            clk_cnt  <= PULSE_WIDTH + HALF_PULSE_WIDTH;
            data_cnt <= 0;
            state    <= STT_DATA;
          end
        end

        default: begin
          state <= STT_WAIT;
        end
      endcase
    end
  end

  assign rx_done = (state == STT_STOP) && (clk_cnt == 0);

  //-----------------------------------------------------------------------------
  // description about output signal



  logic [DATA_WIDTH-1:0] data_r;
  logic                  valid_r;

  always_ff @(posedge clk) begin
    if (!rstn) begin
      data_r  <= 0;
      valid_r <= 0;
    end else if (rx_done && !valid_r) begin
      valid_r <= 1;
      data_r  <= data_tmp_r;
    end else if (valid_r && ready) begin
      valid_r <= 0;
    end
  end

  assign data  = data_r;
  assign valid = valid_r;

endmodule
